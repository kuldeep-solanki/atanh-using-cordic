`timescale 1ns / 1ps

module FloatingDivision(input [31:0]A,input [31:0]B,output [31:0] result);
                         
reg [23:0] A_Mantissa,B_Mantissa;
reg [22:0] Mantissa;
wire [7:0] exp;
reg [23:0] Temp_Mantissa;
reg [7:0] A_Exponent,B_Exponent,Temp_Exponent,diff_Exponent;
wire [7:0] Exponent;
reg [7:0] A_adjust,B_adjust;
reg A_sign,B_sign,Sign;
reg [32:0] Temp;
wire [31:0] temp1,temp2,temp3,temp4,temp5,temp6,temp7,debug;
wire [31:0] reciprocal;
wire [31:0] x0,x1,x2,x3;
reg [6:0] exp_adjust;
reg [31:0] B_scaled; 
reg en1,en2,en3,en4,en5;
reg dummy;
/*----Initial value----*/
FloatingMultiplication M1(.A({{1'b0,8'd126,B[22:0]}}),.B(32'h3ff0f0f1),.result(temp1)); //verified
assign debug = {1'b1,temp1[30:0]};
FloatingAddition A1(32'h4034b4b5,{1'b1,temp1[30:0]},x0);





















/*----First Iteration----*/
FloatingMultiplication M2(.A({{1'b0,8'd126,B[22:0]}}),.B(x0),.result(temp2));
FloatingAddition A2(32'h40000000,{!temp2[31],temp2[30:0]},temp3);
FloatingMultiplication M3(.A(x0),.B(temp3),.result(x1));

/*----Second Iteration----*/
FloatingMultiplication M4(.A({1'b0,8'd126,B[22:0]}),.B(x1),.result(temp4));
FloatingAddition A3(32'h40000000,{!temp4[31],temp4[30:0]},temp5);
FloatingMultiplication M5(.A(x1),.B(temp5),.result(x2));

/*----Third Iteration----*/
FloatingMultiplication M6(.A({1'b0,8'd126,B[22:0]}),.B(x2),.result(temp6));
FloatingAddition A4(32'h40000000,{!temp6[31],temp6[30:0]},temp7);
FloatingMultiplication M7(.A(x2),.B(temp7),.result(x3));

/*----Reciprocal : 1/B----*/
assign Exponent = x3[30:23]+8'd126-B[30:23];
assign reciprocal = {B[31],Exponent,x3[22:0]};

/*----Multiplication A*1/B----*/
FloatingMultiplication M8(.A(A),.B(reciprocal),.result(result));
endmodule



//`timescale 1ns / 1ps

//module FloatingDivision#(parameter XLEN=32)
//                        (input [XLEN-1:0]A,
//                         input [XLEN-1:0]B,
//                         output [XLEN-1:0] result);
                         
//reg [23:0] A_Mantissa,B_Mantissa;
//reg [22:0] Mantissa;
//wire [7:0] exp;
//reg [23:0] Temp_Mantissa;
//reg [7:0] A_Exponent,B_Exponent,Temp_Exponent,diff_Exponent;
//wire [7:0] Exponent;
//reg [7:0] A_adjust,B_adjust;
//reg A_sign,B_sign,Sign;
//reg [32:0] Temp;
//wire [31:0] temp1,temp2,temp3,temp4,temp5,temp6,temp7,debug;
//wire [31:0] reciprocal;
//wire [31:0] x0,x1,x2,x3;
//reg [6:0] exp_adjust;
//reg [XLEN-1:0] B_scaled; 
//reg en1,en2,en3,en4,en5;
//reg dummy;
///*----Initial value----*/
//FloatingMultiplication M1(.A({{1'b0,8'd126,B[22:0]}}),.B(32'h3ff0f0f1),.result(temp1)); //verified
//assign debug = {1'b1,temp1[30:0]};
//FloatingAddition A1(32'h4034b4b5,{1'b1,temp1[30:0]},x0);

///*----First Iteration----*/
//FloatingMultiplication M2(.A({{1'b0,8'd126,B[22:0]}}),.B(x0),.result(temp2));
//FloatingAddition A2(32'h40000000,{!temp2[31],temp2[30:0]},temp3);
//FloatingMultiplication M3(.A(x0),.B(temp3),.result(x1));

///*----Second Iteration----*/
//FloatingMultiplication M4(.A({1'b0,8'd126,B[22:0]}),.B(x1),.result(temp4));
//FloatingAddition A3(32'h40000000,{!temp4[31],temp4[30:0]},temp5);
//FloatingMultiplication M5(.A(x1),.B(temp5),.result(x2));

///*----Third Iteration----*/
//FloatingMultiplication M6(.A({1'b0,8'd126,B[22:0]}),.B(x2),.result(temp6));
//FloatingAddition A4(32'h40000000,{!temp6[31],temp6[30:0]},temp7);
//FloatingMultiplication M7(.A(x2),.B(temp7),.result(x3));

///*----Reciprocal : 1/B----*/
//assign Exponent = x3[30:23]+8'd126-B[30:23];
//assign reciprocal = {B[31],Exponent,x3[22:0]};

///*----Multiplication A*1/B----*/
//FloatingMultiplication M8(.A(A),.B(reciprocal),.result(result));
//endmodule

